

*IDVD
.model MOS NMOS(LEVEL=3 L=2e-06 W=2.3e-05 RSH=30 RS=0.01 RD=0.01 CJ=0 CJSW=0 MJSW=0.33 JS=0 TOX=2e-08 VTO=0.7 PHI=1 GAMMA=1 ETA=0.1 XJ=1e-07 UO=400 THETA=0.001 VMAX=100000 KAPPA=0)

VD D 0 DC 0

VG G 0 DC 0

M1 D G 0 0 MOS

.dc VD 0.0 7.0 0.1 VG LIST 0.4 1.0 1.6 2.2 2.8 3.4 4.0 4.6 5.2 5.8 6.4 7.0
.option plotwinsize=0
.options noopiter

.end

